{"obj/api/nuitrack.PlatformChanger.EnviromentSwitcher.yml":{"~/obj/api/nuitrack.PlatformChanger.EnviromentSwitcher.yml":"~/api/nuitrack.PlatformChanger.EnviromentSwitcher.html"},"obj/api/nuitrack.Pointer.PointerPassing.CalibrationAction.yml":{"~/obj/api/nuitrack.Pointer.PointerPassing.CalibrationAction.yml":"~/api/nuitrack.Pointer.PointerPassing.CalibrationAction.html"},"obj/api/nuitrack.VicoVRCalibration.yml":{"~/obj/api/nuitrack.VicoVRCalibration.yml":"~/api/nuitrack.VicoVRCalibration.html"},"obj/api/nuitrack.Frame.DepthToTexture.yml":{"~/obj/api/nuitrack.Frame.DepthToTexture.yml":"~/api/nuitrack.Frame.DepthToTexture.html"},"obj/api/User.yml":{"~/obj/api/User.yml":"~/api/User.html"},"obj/api/nuitrack.Frame.yml":{"~/obj/api/nuitrack.Frame.yml":"~/api/nuitrack.Frame.html"},"obj/api/nuitrack.Pointer.yml":{"~/obj/api/nuitrack.Pointer.yml":"~/api/nuitrack.Pointer.html"},"obj/api/nuitrack.VicoVRCalibration.SensorDisconnectChecker.yml":{"~/obj/api/nuitrack.VicoVRCalibration.SensorDisconnectChecker.yml":"~/api/nuitrack.VicoVRCalibration.SensorDisconnectChecker.html"},"obj/api/nuitrack.PlatformChanger.GameVersion.yml":{"~/obj/api/nuitrack.PlatformChanger.GameVersion.yml":"~/api/nuitrack.PlatformChanger.GameVersion.html"},"obj/api/nuitrack.Pointer.PointerPassing.ClickAction.yml":{"~/obj/api/nuitrack.Pointer.PointerPassing.ClickAction.yml":"~/api/nuitrack.Pointer.PointerPassing.ClickAction.html"},"obj/api/nuitrack.VicoVRCalibration.SensorDisconnectChecker.ConnectionStatusChange.yml":{"~/obj/api/nuitrack.VicoVRCalibration.SensorDisconnectChecker.ConnectionStatusChange.yml":"~/api/nuitrack.VicoVRCalibration.SensorDisconnectChecker.ConnectionStatusChange.html"},"obj/api/nuitrack.Frame.SegmentToTexture.yml":{"~/obj/api/nuitrack.Frame.SegmentToTexture.yml":"~/api/nuitrack.Frame.SegmentToTexture.html"},"obj/api/nuitrack.Pointer.PointerPassing.yml":{"~/obj/api/nuitrack.Pointer.PointerPassing.yml":"~/api/nuitrack.Pointer.PointerPassing.html"},"obj/api/nuitrack.VicoVRCalibration.BackTextureCreator.yml":{"~/obj/api/nuitrack.VicoVRCalibration.BackTextureCreator.yml":"~/api/nuitrack.VicoVRCalibration.BackTextureCreator.html"},"obj/api/nuitrack.Frame.TextureCache.yml":{"~/obj/api/nuitrack.Frame.TextureCache.yml":"~/api/nuitrack.Frame.TextureCache.html"},"obj/api/nuitrack.Pointer.PointerRotation.yml":{"~/obj/api/nuitrack.Pointer.PointerRotation.yml":"~/api/nuitrack.Pointer.PointerRotation.html"},"obj/api/User.UserAvatar.yml":{"~/obj/api/User.UserAvatar.yml":"~/api/User.UserAvatar.html"},"obj/api/nuitrack.Frame.FrameOverloadUtils.yml":{"~/obj/api/nuitrack.Frame.FrameOverloadUtils.yml":"~/api/nuitrack.Frame.FrameOverloadUtils.html"},"obj/api/nuitrack.VicoVRCalibration.BackTextureCreator.newBackGroundCreate.yml":{"~/obj/api/nuitrack.VicoVRCalibration.BackTextureCreator.newBackGroundCreate.yml":"~/api/nuitrack.VicoVRCalibration.BackTextureCreator.newBackGroundCreate.html"},"obj/api/User.UserAvatar.Connection.yml":{"~/obj/api/User.UserAvatar.Connection.yml":"~/api/User.UserAvatar.Connection.html"},"obj/api/nuitrack.Frame.FrameUtils.yml":{"~/obj/api/nuitrack.Frame.FrameUtils.yml":"~/api/nuitrack.Frame.FrameUtils.html"},"obj/api/nuitrack.Pointer.VVRInput.yml":{"~/obj/api/nuitrack.Pointer.VVRInput.yml":"~/api/nuitrack.Pointer.VVRInput.html"},"obj/api/nuitrack.VicoVRCalibration.RGBCalibrationVisualizer.yml":{"~/obj/api/nuitrack.VicoVRCalibration.RGBCalibrationVisualizer.yml":"~/api/nuitrack.VicoVRCalibration.RGBCalibrationVisualizer.html"},"obj/api/nuitrack.Frame.FrameToTexture-2.yml":{"~/obj/api/nuitrack.Frame.FrameToTexture-2.yml":"~/api/nuitrack.Frame.FrameToTexture-2.html"},"obj/api/nuitrack.Pointer.VVRInput.Button.yml":{"~/obj/api/nuitrack.Pointer.VVRInput.Button.yml":"~/api/nuitrack.Pointer.VVRInput.Button.html"},"obj/api/Ray.yml":{"~/obj/api/Ray.yml":"~/api/Ray.html"},"obj/api/nuitrack.PlatformChanger.yml":{"~/obj/api/nuitrack.PlatformChanger.yml":"~/api/nuitrack.PlatformChanger.html"},"obj/api/nuitrack.SafetyGrid.SensorPointReplacer.yml":{"~/obj/api/nuitrack.SafetyGrid.SensorPointReplacer.yml":"~/api/nuitrack.SafetyGrid.SensorPointReplacer.html"},"obj/api/nuitrack.Frame.RGBToTexture.yml":{"~/obj/api/nuitrack.Frame.RGBToTexture.yml":"~/api/nuitrack.Frame.RGBToTexture.html"},"obj/api/nuitrack.SafetyGrid.yml":{"~/obj/api/nuitrack.SafetyGrid.yml":"~/api/nuitrack.SafetyGrid.html"},"obj/api/Ray.RayScript.yml":{"~/obj/api/Ray.RayScript.yml":"~/api/Ray.RayScript.html"},"obj/api/nuitrack.Frame.TextureUtils.yml":{"~/obj/api/nuitrack.Frame.TextureUtils.yml":"~/api/nuitrack.Frame.TextureUtils.html"},"obj/api/nuitrack.Pointer.PointerVisuals.yml":{"~/obj/api/nuitrack.Pointer.PointerVisuals.yml":"~/api/nuitrack.Pointer.PointerVisuals.html"},"index.md":{"~/index.md":"~/index.html"},"api/index.md":{"~/api/index.md":"~/api/index.html"},"articles/intro.md":{"~/articles/intro.md":"~/articles/intro.html"},"articles/toc.md":{"~/articles/toc.md":"~/articles/toc.html"},"toc.yml":{"~/toc.yml":"~/toc.html"},"obj/api/toc.yml":{"~/obj/api/toc.yml":"~/api/toc.html"}}